`include "def.h"

module stack(clk, reset, load, push, pop, d, qtop, qnext);

    
