`include "def.h"

module alu(
input [`DATA_W-1:0] a,b,
input [`OPCODE_W-1:0] s,
output [`DATA_W-1:0] o);

endmodule
